---- The Data Path
--
--library ieee;
--
--use ieee.std_logic_arith.all;
--use ieee.std_logic_1164.all;
--
--
--Entity datapath is
--    Port(clk        : in std_logic;
--         reset      : in std_logic;
--         memtoreg   : in std_logic;
--         pcsrc      : in std_logic;
--         alusrc     : in std_logic;
--         regdst     : in std_logic;
--         regwrite   : in std_logic;
--         alucontrol : in std_logic_vector(3 downto 0);
--         instruction: in std_logic_vector(31 downto 0);
--         readdata   : in std_logic_vector(31 downto 0);
--         pc         : out std_logic_vector(31 downto 0);
--         aluout     : out std_logic_vector(31 downto 0);
--         writedata  : out std_logic_vector(31 downto 0);
--         zero       : out std_logic);
--end datapath;
--
--architecture behaviour of datapath is
--
--    component ControlUnit
--	port(opcode : in std_logic_vector (5 DOWNTO 0);
--		ALUOp : out std_logic_vector(5 DOWNTO 0);
--		regDst, memRead, memToRegister, memWrite, ALUsrc, regWrite : out std_logic);
--	end component;
--	for ctrlUnit: ControlUnit use entity work.ControlUnit;
--
--    component alu
--    port(a1       : in std_logic_vector(31 downto 0);
--         a2       : in std_logic_vector(31 downto 0);
--         alu_control : in std_logic_vector(3 downto 0);
--         alu_result  : out std_logic_vector(31 downto 0);
--         zero       : out std_logic);
--    end component;
--    for alu0: alu use entity work.alu;
--
--    component alu_control
--	port(ALUOp : in STD_LOGIC_VECTOR (5 DOWNTO 0);
--	     operation : OUT std_logic_vector (3 DOWNTO 0));
--    end component;
--    for aluCtrl: alu_control use entity work.alu_control;
--
--    component REGISTER_FILE
--        port(readRegister1  : in std_logic_vector(4 downto 0);
--            readRegister2  : in std_logic_vector(4 downto 0);
--	    readData1 : out std_logic_vector(31 downto 0);
--            readData2 : out std_logic_vector(31 downto 0);
--	     registerWrite : in std_logic;
--            writeData : in std_logic_vector(31 downto 0));
--            --clk : in std_logic; may add
--            
--    end component;
--    for rf0 : REGISTER_FILE use entity work.REGISTER_FILE;
--
--    component PC_ADDER
--        port(PC_IN : in std_logic_vector(31 downto 0);
--             PC_OUT    : out std_logic_vector(31 downto 0));
--    end component;
--    for pcadder : adder use entity work.PC_ADDER;
--
--    component SIGN_EXTENDER
--        port(numIn : in std_logic_vector(15 downto 0);
--             numOut : out std_logic_vector(31 downto 0));
--    end component;
--    for signext0 : SIGN_EXTENDER use entity work.SIGN_EXTENDER;
--
--    component TwoToOneMux;
--        port(in0, in1 : in std_logic_vector(31 downto 0);
--             out0      : out std_logic_vector(31 downto 0);
--	     cSwitch      : in std_logic);
--    end component;
--    for muxregdest : mux use entity work.mux;
--    for muxalusrc : mux use entity work.mux;
--    for muxaluout : mux use entity work.mux;
--
--    component IFToID
--    Port (clk         : in std_logic;
--	  instruction : in std_logic_vector(31 downto 0);
--	  OpCode      : out std_logic(5 downto 0);
--	  readRegister1 : out std_logic_vector(4 downto 0);
--	  readRegister2 : out std_logic_vector(4 downto 0);
--          immediateValue : out std_logic_vector(4 downto 0);
--	  IwriteRegister : out std_logic_vector(4 downto 0);
--	  RwriteRegister : out std_logic_vector(4 downto 0));
--    end component;
--    for regpipe1 : IFToID use entity work.IDToID;
--
--    component IDToEX 
--    Port (clk : IN std_logic;
--		-- Inputs
--				
--		ALUopIN	      	  : IN std_logic_vector(5 DOWNTO 0); -- same as opcode
--		regDstIN          : IN std_logic; -- 0 for immediate and LW/SW, 1 for register arith
--		memReadIN         : IN std_logic; -- 1 for reading memory
--		memToRegisterIN   : IN std_logic; -- 1 for memRead data goes to destination register else 0 for ALU result to destination register
--		memWriteIN        : IN std_logic; -- 1 for writing data
--		ALUsrcIN          : IN std_logic; -- 0 for second operand to be a register else 1 for second operand is immediate value (direct value offest for a mem address)
--		regWriteIN  	  : IN std_logic;  -- 1 for computed result is written to destination register, in this project only 0 for SW
--		readData1IN       : IN std_logic_vector (31 DOWNTO 0);-- Data read from register 1
--		readData2IN       : IN std_logic_vector (31 DOWNTO 0);-- Data read from register 2
--		signExtendIN  	  : IN STD_logic_vector(31 DOWNTO 0);  -- the extended number
--		IwriteRegisterIN  : IN std_logic_vector (4 DOWNTO 0);  -- Register where where data will be written to if "I" instruction
--		RwriteRegisterIN  : IN std_logic_vector (4 DOWNTO 0);  -- Register where where data will be written to if "R" instruction
--
--		-- Outputs (same as Inputs)
--		ALUopOUT	   : OUT std_logic_vector(5 DOWNTO 0); -- same as opcode
--		regDstOUT          : OUT std_logic; -- 0 for immediate and LW/SW, 1 for register arith
--		memReadOUT         : OUT std_logic; -- 1 for reading memory
--		memToRegisterOUT   : OUT std_logic; -- 1 for memRead data goes to destination register else 0 for ALU result to destination register
--		memWriteOUT        : OUT std_logic; -- 1 for writing data
--		ALUsrcOUT          : OUT std_logic; -- 0 for second operand to be a register else 1 for second operand is immediate value (direct value offest for a mem address)
--		regWriteOUT  	   : OUT std_logic;  -- 1 for computed result is written to destination register, in this project only 0 for SW
--		readData1OUT       : OUT std_logic_vector (31 DOWNTO 0);-- Data read from register 1
--		readData2OUT       : OUT std_logic_vector (31 DOWNTO 0);-- Data read from register 2
--		signExtendOUT  	   : OUT STD_logic_vector(31 DOWNTO 0);  -- the extended number
--		IwriteRegisterOUT  : OUT std_logic_vector (4 DOWNTO 0);  -- Register where where data will be written to if "I" instruction
--		RwriteRegisterOUT  : OUT std_logic_vector (4 DOWNTO 0)  -- Register where where data will be written to if "R" instruction
--		
--	);
--    end component;
--    for regpipe2 : IDToEx use entity work.IDToEX;
--
--    component EXToMEM
--    Port (clk : IN std_logic;
--		-- Input
--		memReadIN         : IN std_logic; -- 1 for reading memory
--		memToRegisterIN   : IN std_logic; -- 1 for memRead data goes to destination register else 0 for ALU result to destination register
--		memWriteIN        : IN std_logic; -- 1 for writing data
--		regWriteIN  	  : IN std_logic;  -- 1 for computed result is written to destination register, in this project only 0 for SW
--		readData2IN       : IN std_logic_vector (31 DOWNTO 0);-- Data read from register 
--		ALUResultIN 	  : IN std_logic_vector (31 DOWNTO 0);-- Computed result from ALU
--		writeRegisterIN   : IN std_logic_vector (4 DOWNTO 0);  -- Register where where data will be written to (Came from multiplexer between IwriteRegister and RwriteRegister)
--
--		-- Outputs (same as Inputs)
--		memReadOUT         : OUT std_logic; -- 1 for reading memory
--		memToRegisterOUT   : OUT std_logic; -- 1 for memRead data goes to destination register else 0 for ALU result to destination register
--		memWriteOUT        : OUT std_logic; -- 1 for writing data
--		regWriteOUT  	   : OUT std_logic;  -- 1 for computed result is written to destination register, in this project only 0 for SW
--		readData2OUT       : OUT std_logic_vector (31 DOWNTO 0);-- Data read from register 2
--		ALUResultOUT 	   : OUT std_logic_vector (31 DOWNTO 0);-- Computed result from ALU
--		writeRegisterOUT   : OUT std_logic_vector (4 DOWNTO 0)  -- Register where where data will be written to (Came from multiplexer between IwriteRegister and RwriteRegister)
--		
--	);
--    end component;
--    for regpipe3 : EXToMEM use entity work.EXToMEM;
--
--    component MEMToWB
--    Port (clk : IN std_logic;
--		-- Inputs
--				
--		memToRegisterIN   : IN std_logic; -- 1 for memRead data goes to destination register else 0 for ALU result to destination register
--		regWriteIN  	  : IN std_logic;  -- 1 for computed result is written to destination register, in this project only 0 for SW
--		readData2IN       : IN std_logic_vector (31 DOWNTO 0);-- Data read from register 2 (it is the write data)
--		ALUResultIN 	  : IN std_logic_vector (31 DOWNTO 0);-- Computed result from ALU
--		writeRegisterIN   : IN std_logic_vector (4 DOWNTO 0);  -- Register where where data will be written to (Came from multiplexer between IwriteRegister and RwriteRegister)
--
--		-- Outputs (same as Inputs)
--		
--		memToRegisterOUT   : OUT std_logic; -- 1 for memRead data goes to destination register else 0 for ALU result to destination register
--		regWriteOUT  	   : OUT std_logic;  -- 1 for computed result is written to destination register, in this project only 0 for SW
--		readData2OUT       : OUT std_logic_vector (31 DOWNTO 0);-- Data read from register 2 (it is the write data)
--		ALUResultOUT 	   : OUT std_logic_vector (31 DOWNTO 0);-- Computed result from ALU
--		writeRegisterOUT   : OUT std_logic_vector (4 DOWNTO 0)  -- Register where where data will be written to (Came from multiplexer between IwriteRegister and RwriteRegister)
--		
--	);
--    end component;
--    for regpipe4 : MEMToWB use entity work.MEMToWB;
--
--    Component PROGRAM_COUNTER
--    Port (clk : in std_logic;
--          PC_IN   : in std_logic_vector(31 downto 0);
--          PC_OUT   : out std_logic_vector(31 downto 0));
--    end component;
--    for pcreg : PROGRAM_COUNTER use entity work.PROGRAM_COUNTER;
--
---- edit these signals
--    signal writereg, writerege, writeregm, writeregW  : std_logic_vector(4 downto 0);
--    signal instructiond, instructionE, ReadDataW, writedataE, writedM : std_logic_vector(31 downto 0);
--    signal memtoregE, memtoregM, memtoregW, alusrcE, memwrite : std_logic;
--    signal ZeroE, regwriteE, regwriteM, regwriteW, regdstE : std_logic;
--    signal alucontrolE : std_logic_vector(2 downto 0);
--    signal pcjump, pcnext, pcnextbr, pcbranchE, pcbranchM, sigimnE, srcae,
--           pcplus4, pcbranch, sigimn, aluoutM, aluoutW, pcplus4D, pcplus4E,
--           signimsh, srca, srcb, result : std_logic_vector(31 downto 0);
--    signal temp : std_logic_vector(31 downto 0);
--
--    signal 
--
--    begin
--        -- IF
--  
--        pcreg : program_counter port map(clk, pcnext, temp); -- pc 
--        pc <= temp; 
--        pcadder : pc_adder port map(temp, pcplus4); -- 
--        regpipe1 : IFToID port map(clk, instruction -- assign signals to outputs);
--
--        -- ID
--
--        rf0 : REGISTER_FILE port map(instructionD(25 downto 21), instructionD(20 downto 16), srca, temp, regwrite, writereg, result); -- Register File
--        writedata <= temp;
--        signext0: signextension port map(instructionD(15 downto 0), sigimn); -- extende imediato
--        regpipe2 : IDToEX port map(clk, regwrite, memtoreg, memwrite, pcbranch, alucontrol, alusrc, regdst, srca, temp,
--                                    instructionD(20 downto 16), instructionD(15 downto 11), sigimn, pcplus4D,
--                                    regwriteE, memtoregE, memwrite, pcbranchE, alucontrolE, alusrcE, regdstE, srcaE, writedataE, 
--                                    instructionD(20 downto 16), instructionE(15 downto 11), sigimnE, pcplus4E);
--
--        -- EX
--
--        muxalusrc: mux generic map(32) port map(writedataE, sigimnE, alusrcE, srcb); -- qual entrada de scrb da alu
--        muxregdest:mux generic map(5) port map(instructionE(20 downto 16), instructionE(15 downto 11), regdstE, writereg);
--        alu0 : alu port map(srca, srcb, alucontrolE, aluout, zeroE); -- verificar se nao precisa de caryout e valores
--        aluout <= temp;
--        regpipe3 : regaux3 generic map(32) port map(clk, regwriteE, memtoregE, memwrite, pcbranchE, zeroE, temp, writedatae, writereg, pcbranchE,
--                                        regwriteM, memtoregM, memwrite, pcbranchM, zero, aluoutM, writedM, writeregM, pcbranchM);
--
--        -- MEM
--
--        regpipe4 : regaux4 generic map(32) port map(clk, regwriteM, memtoregM, readdata, aluoutM, writeregM, regwriteW, memtoregW, readdataW, aluoutW, writeregW);
--        -- WB
--
--        muxaluout : mux generic map(32) port map(readdataW, aluoutW, memtoregW, result);
--
--
--end behaviour;
